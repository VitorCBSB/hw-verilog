module sender();

	

endmodule